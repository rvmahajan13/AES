library ieee;
use ieee.std_logic_1164.all;

package Utilities is 
	type matrix is array(0 to 3, 0 to 3) of std_logic_vector(7 downto 0);
end package;